module test_lena;

tester tester();

endmodule

