module test_image3;

tester tester();

endmodule

