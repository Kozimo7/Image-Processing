module test_image2;

tester tester();

endmodule

